  module memory (dout, insn, addr, insn_addr, clk, din, mem_we);

	//read_addr and write_addr combined
	input [31:0] insn_addr, addr, din;
	input [3:0] mem_we;
	input clk;
	output reg [31:0] dout, insn;

	reg [31:0] mem [0:1023]; //Little Endian

	/*INITIALISATION

	initial 
		begin
	    	for (i=0; i < 1024; i=i+1) 
	    		begin
		 			mem[i] = 32'b0;
	      		end

		mem[0] = 32'b00000000000100000000001010010011;
		mem[1] = 32'b00000000000100101000001010010011;
		mem[2] = 32'b00000000001100000000001010010011;
		mem[3] = 32'b00000000000100101000001010010011;
		mem[4] = 32'b11111111111100000000001010010011;
		mem[5] = 32'b00000000000100101000001010010011;
		mem[6] = 32'b00000000000100000000000000010011;
		mem[7] = 32'b00000000000100000000000010010011;
		mem[8] = 32'b00000000000100001000000100010011;
		mem[9] = 32'b00000000000100010000000110010011;
		mem[10] = 32'b00000000000100011000001000010011;
		mem[11] = 32'b00000000000100100000001010010011;
		mem[12] = 32'b00000000000100101000001100010011;
		mem[13] = 32'b00000000000100110000001110010011;
		mem[14] = 32'b00000000000100111000010000010011;
		mem[15] = 32'b00000000000101000000010010010011;
		mem[16] = 32'b00000000000101001000010100010011;
		mem[17] = 32'b00000000000101010000010110010011;
		mem[18] = 32'b00000000000101011000011000010011;
		mem[19] = 32'b00000000000101100000011010010011;
		mem[20] = 32'b00000000000101101000011100010011;
		mem[21] = 32'b00000000000101110000011110010011;
		mem[22] = 32'b00000000000101111000100000010011;
		mem[23] = 32'b00000000000110000000100010010011;
		mem[24] = 32'b00000000000110001000100100010011;
		mem[25] = 32'b00000000000110010000100110010011;
		mem[26] = 32'b00000000000110011000101000010011;
		mem[27] = 32'b00000000000110100000101010010011;
		mem[28] = 32'b00000000000110101000101100010011;
		mem[29] = 32'b00000000000110110000101110010011;
		mem[30] = 32'b00000000000110111000110000010011;
		mem[31] = 32'b00000000000111000000110010010011;
		mem[32] = 32'b00000000000111001000110100010011;
		mem[33] = 32'b00000000000111010000110110010011;
		mem[34] = 32'b00000000000111011000111000010011;
		mem[35] = 32'b00000000000111100000111010010011;
		mem[36] = 32'b00000000000111101000111100010011;
		mem[37] = 32'b00000000000111110000111110010011;
		mem[38] = 32'b00000000000000000000000001101111;
	      
	    end

    */

	always @(posedge clk) 
		begin
			if(clk&mem_we)
				begin
					//mem[addr]<=din; addr[9:0] because 2^10=1024
					mem[addr[11:2]][7:0] <= mem_we[0] ? din[7:0] : mem[addr[9:0]][7:0];
      				mem[addr[11:2]][15:8] <= mem_we[1] ? din[15:8] : mem[addr[9:0]][15:8];
      				mem[addr[11:2]][23:16] <= mem_we[2] ? din[23:16] : mem[addr[9:0]][23:16];
      				mem[addr[11:2]][31:24] <= mem_we[3] ? din[31:24] : mem[addr[9:0]][31:24];
				end
			dout = mem[addr[11:2]];
			insn = mem[insn_addr[11:2]];
		end       

endmodule
